parameter tag_length = 5;
parameter addr_width = 8;
parameter data_width = 32;

typedef enum bit {RD,WR} tx_type_e;
