typedef uvm_sequencer#(axi_seq_item) axi_sqr;
